-- Testbench for logic gates
