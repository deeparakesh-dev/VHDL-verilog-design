-- Logic gates design 
