-- Logic gates design 
--AND,OR,NOT,XOR,XNOR,NAND
